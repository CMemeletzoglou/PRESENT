LIBRARY ieee;
USE ieee.std_logic_1164.all;

package key_length_pack is
        -- type KEY_LENGTH is (KEY_80, KEY_128);
        constant KEY_LENGTH : NATURAL := 80;        
end package;