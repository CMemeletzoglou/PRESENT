LIBRARY ieee;
USE ieee.std_logic_1164.all;

package key_length_pkg is
--        constant KEY_LENGTH : NATURAL := 80;
       constant KEY_LENGTH : NATURAL := 128;
end package;