library ieee;
use ieee.std_logic_1164.all;

entity present_enc is
        port (
                clk               : in std_logic;
                rst               : in std_logic;
                ena               : in std_logic;
                plaintext         : in std_logic_vector(63 downto 0);
                round_key         : in std_logic_vector(63 downto 0); -- read from round keys mem
                current_round_num : out std_logic_vector(4 downto 0);
                ciphertext        : out std_logic_vector(63 downto 0);
                ready             : out std_logic
        );
end present_enc;

architecture structural of present_enc is
        constant BLOCK_SIZE : natural := 64;

        signal  mux_sel,
                ciph_enable : std_logic;

        signal  state_reg_mux_out,
                state : std_logic_vector(BLOCK_SIZE - 1 downto 0);

        signal  sbox_layer_input,
                pbox_layer_input,
                pbox_layer_out : std_logic_vector(BLOCK_SIZE - 1 downto 0);

        signal  key_reg_out : std_logic_vector(BLOCK_SIZE - 1 downto 0);

        signal  round_num : std_logic_vector(4 downto 0);
begin
        -- control signal for the multiplexers controlling the input of
        -- State and Key registers
        mux_sel <= '1' when (round_num = "00000") else '0';

        -- 64-bit mux which drives the state register
        state_reg_mux : entity work.mux
                generic map(
                        DATA_WIDTH => BLOCK_SIZE
                )
                port map(
                        input_A => pbox_layer_out,
                        input_B => plaintext,
                        sel     => mux_sel,
                        mux_out => state_reg_mux_out
                );

        -- 64-bit state register
        state_reg : entity work.reg
                generic map(
                        DATA_WIDTH => BLOCK_SIZE
                )
                port map(
                        clk  => clk,
                        rst  => rst,
                        ena  => ena,
                        din  => state_reg_mux_out,
                        dout => state
                );

        -- 64-bit key register, it stores the current round key retrieved from the round keys memory
        -- TODO : unecessary (??)
        key_reg : entity work.reg
                generic map(
                        DATA_WIDTH => 64
                )
                port map(
                        clk  => clk,
                        rst  => rst,
                        ena  => ena,
                        din  => round_key,
                        dout => key_reg_out
                );

        -- 64-bit xor to add current round key to state
        xor_64 : entity work.xor_n
                generic map(
                        DATA_WIDTH => BLOCK_SIZE
                )
                port map(
                        a => state,
                        b => key_reg_out,
                        y => sbox_layer_input
                );

        -- S-Box layer (16 S-Boxes in parallel), the *confusion* layer
        sbox_layer : entity work.sbox_layer
                port map(
                        sbox_layer_in  => sbox_layer_input,
                        sbox_layer_out => pbox_layer_input
                );

        -- P-Box layer, the *diffusion* layer
        pbox_layer : entity work.pbox
                port map(
                        data_in  => pbox_layer_input,
                        data_out => pbox_layer_out
                );

        -- round counter, incremented by 1 at each network round
        round_counter : entity work.counter
                generic map(
                        COUNTER_WIDTH => 5
                )
                port map(
                        clk    => clk,
                        rst    => rst,
                        ena    => ena,
                        updown => '0',
                        count  => round_num
                );

        current_round_num <= round_num;

        -- 64-bit ciphertext register
        ciph_reg : entity work.reg
                generic map(
                        DATA_WIDTH => BLOCK_SIZE
                )
                port map(
                        clk  => clk,
                        rst  => rst,
                        ena  => ciph_enable,
                        din  => sbox_layer_input,
                        dout => ciphertext
                );

        -- ciphertext register enable signal, must be activated when the
        -- round_counter overflows to "00000". Since the output of the
        -- round_counter is a signal, the value read from it is one cycle behind.
        -- So the round_counter is found to be "00000", during the first round of
        -- the next encryption cycle. So we need 31 cycles for the actual encryption
        -- + 1 cycle to get the encrypted plaintext on the ciphertext output bus
        with round_num select
                ciph_enable <= '1' when "00000",
                '0' when others;

        -- when round_counter overflows to "00000", we are finished
        -- so raise the finished flag, indicating that the contents of
        -- the ciphertext output are valid and correspond to the 
        -- encrypted plaintext. Compare the round_counter to "00001" and not to
        -- "00000" as in the select statement above, in order to give the ciphertext
        -- register, the necessary cycle to pass the ciphertext from its input to its 
        -- output
        with round_num select
                ready <= '1' when "00001",
                '0' when others;

        -- small issue though.. the ready flag is also raised during the first encryption
        -- process' second cycle (counter = 000001)
end structural;