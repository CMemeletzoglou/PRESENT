package state_pkg is
        type STATE is (INIT, KEY_GEN, CRYPTO_OP, DONE, INVALID);
end package;
